
module addbit (
a, 
b, 
cin, 
sum, 
cout
);


input a;
input b;
input cin;
output sum;
output cout;

assign {co,sum} = a + b + ci;

endmodule
